`define BUS 31:0
`define BUSW 32
`define BUSWT 31 
`define BUS_REG 4:0
`define BUS_ADDR 23:0
`define BUS_ADDRW 24
`define BUS_ADDRWT 23