`define BUS 31:0
`define BUS_REG 4:0