`define BUS 31:0
`define BUSW 32
`define BUSWT 31 
`define BUS_REG 4:0